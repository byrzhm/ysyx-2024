module ysyx_22040000_IFU (
    input [31:0] pc,
    output reg [31:0] inst
);

    // TODO

endmodule
